library ieee;
use ieee.std_logic_1164.all;


package Pack is

	type instruction_type is (DP_R, DP_I, LS, BBL, S);

end Pack;


